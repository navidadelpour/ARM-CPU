module PcTestbench ();

	ALU(